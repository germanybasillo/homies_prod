b0VIM 8.2      �ag)+ G  Administrator                           PC01                                    /c/laragon/www/lagotlagot/resources/views/welcome.blade.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           W                            $       X                     F       }                     h       �                     Z       *                    g       �             	       V       �             
       m       A                    X       �                    Q                           f       W                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     �     W       �  �  N    �  �  �  �  �  =  *  �  �  �  �  `  N  �  �  �  k  ]    �  |    �
  �
  ]
  !
  
  �	  �	  �	  o	  -	  	  �  �  }    �  �  �  �  �  {  T  5  �  �  �  �  �  �  i  W  ,  �  �  �  Y    �  �  �  }  s  o  n  N  1  0    �  �  �  �  �  �  �  �  �  L  *     �  �                            <a href="/" class="navbar-brand scroll-top logo  animated bounceInLeft"><b><i><img src="/logo.png" style="height: 60px;"/></i></b></a> </div>         <button type="button" id="nav-toggle" class="navbar-toggle" data-toggle="collapse" data-target="#main-nav"> <span class="sr-only">Toggle navigation</span> <span class="icon-bar"></span> <span class="icon-bar"></span> <span class="icon-bar"></span> </button>       <div class="navbar-header">     <nav class="navbar navbar-inverse" role="navigation">   <div class="container"> <header class="header"> <body>  </head>   </script>   window.addEventListener('offline', showNoInternetMessage);   // Listen for offline events    checkInternetConnection();   // Initial check on page load    }       });           }               location.reload(); // Reload the page on confirmation           if (result.isConfirmed) {       }).then((result) => {           allowEscapeKey: false // Prevents closing by using the escape key           allowOutsideClick: false, // Prevents closing by clicking outside           confirmButtonText: 'Reload',           icon: 'warning',           text: 'Please check your connection and reload the page.',           title: 'No Internet Connection',       Swal.fire({   function showNoInternetMessage() {   // Function to show a "No Internet" message using SweetAlert2    }       }           showNoInternetMessage();           // If no internet connection, show a message       if (!navigator.onLine) {   function checkInternetConnection() {   // Function to check if the browser is offline <script>    <script src="https://unpkg.com/leaflet-control-geocoder/dist/Control.Geocoder.js"></script>  <link rel="stylesheet" href="https://unpkg.com/leaflet-control-geocoder/dist/Control.Geocoder.css" />   crossorigin=""></script>   integrity="sha256-20nQCchB9co0qIjJZRGuk2/Z9VM+kNiyxNV1lvTlZBo="   <script src="https://unpkg.com/leaflet@1.9.4/dist/leaflet.js"   crossorigin=""/>   integrity="sha256-p4NxAoJBhIIN+hmNHrzRCf9tD/miZyoHS5obTRR9BMY="   <link rel="stylesheet" href="https://unpkg.com/leaflet@1.9.4/dist/leaflet.css"     <link href="landingpage/font/css/font-awesome.min.css" rel="stylesheet"> <!-- Font Awesome --> <link rel="stylesheet" href="landingpage/css/styles.css" /> <link href="landingpage/js/owl-carousel/owl.carousel.css" rel="stylesheet"> <!-- Owl Carousel Assets --> <link href="landingpage/css/animate.css" rel="stylesheet" media="screen"> <link rel="stylesheet" href="landingpage/js/fancybox/jquery.fancybox.css" type="text/css" media="screen" /> <link rel="stylesheet" type="text/css" href="landingpage/css/isotope.css" media="screen" /> <link rel="icon" href="{{ asset('logo.png') }}" type="image/png"> <link rel="stylesheet" href="landingpage/css/bootstrap.min.css" /> 	<![endif]--> 		<script type="text/javascript" src="http://explorercanvas.googlecode.com/svn/trunk/excanvas.js"></script> <!--[if lte IE 8]>     <![endif]-->         <script src="http://html5shim.googlecode.com/svn/trunk/html5.js"></script> <!--[if lt IE 9]> <meta name="author" content="WebThemez"> <meta name="description" content=""> <title>{{ config('app.name') }}</title>     <![endif]-->     <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1"> <!--[if lt IE 9]>  <meta name="viewport" content="width=device-width, initial-scale=1, maximum-scale=1"> <meta charset="utf-8"> <head> <!--<![endif]--> <html lang="en-gb" class="no-js"> <!--[if (gt IE 9)|!(IE)]><!--> <!--[if IE 9 ]>    <html lang="en-gb" class="isie ie9 no-js"> <![endif]--> <!--[if IE 8 ]>    <html lang="en-gb" class="isie ie8 oldie no-js"> <![endif]--> <!--[if IE 7 ]>    <html lang="en-gb" class="isie ie7 oldie no-js"> <![endif]--> <!doctype html> ad  R  �            �  �  �  �  �  |  Q    �  �  ~  2    �  �  �  �  �  �  s  V  U  6  �  �  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    </html> </body>  </script>   window.addEventListener('offline', showNoInternetMessage);   // Listen for offline events    checkInternetConnection();   // Initial check on page load    }       });           }               location.reload(); // Reload the page on confirmation           if (result.isConfirmed) {       }).then((result) => {           allowEscapeKey: false // Prevents closing by using the escape key           allowOutsideClick: false, // Prevents closing by clicking outside           confirmButtonText: 'Reload',           icon: 'warning',           text: 'Please check your connection and reload the page.',           title: 'No Internet Connection',       Swal.fire({   function showNoInternetMessage() {   // Function to show a "No Internet" message using SweetAlert2    }       } ad  S  �     F       �  �  o  f  I    �  �  �  �  ?  !    �  �  �  �  �  }  k  [  Z  �  �  s  N  �  �  �  �  �  �  �  �  t  k  U  K  ;  %    �
  �
  {
  4
  �	  �	  �	  �	  �	  v	  1	  �  �  �  �  �  �  f  G  (  	  �  �  �  �  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         @php  @endforeach   @endphp       ]);           $selected->profile6           $selected->profile5,           $selected->profile4,           $selected->profile2,           $selected->profile1,           $selected->profile3,       $images = array_merge($images, [       // Collect all profile images into the array   @php @foreach($selecteds as $selected)  @endphp   $images = []; // Initialize an empty array to collect images   $selecteds = App\Models\Selected::inRandomOrder()->take(3)->get();   // Fetch 3 random selected records   @php   <!-- Carousel items -->   </ol>     <li data-target="#carousel" data-slide-to="2"></li>     <li data-target="#carousel" data-slide-to="1"></li>     <li data-target="#carousel" data-slide-to="0" class="active"></li>   <ol class="carousel-indicators">   	<div id="carousel" class="carousel slide carousel-fade" data-ride="carousel">   <div class="banner-container">  <section id="home"> <div id="#top"></div> <!--/.header--> </header>   <!--/.container-->    </div>     <!--/.navbar-->      </nav>       <!--/.navbar-collapse-->        </div>     </ul>     @endif         @endauth         @endif             <li><a href="{{ route('register') }}" class="scroll-link">Register</a></li>         @if (Route::has('register'))         <li><a href="{{ route('login') }}" class="scroll-link">Login</a></li>     @else         <li><a href="#" onclick="event.preventDefault(); document.getElementById('logout-form').submit();" class="scroll-link">Logout</a></li>          </form>             @csrf         <form id="logout-form" action="{{ route('logout') }}" method="POST" style="display: none;">  </script>     });         }             });                 );                     'warning'                     'Your account is still pending. Please wait for approval.',                     'Account Pending',                 Swal.fire(                                  e.preventDefault();             dashboardLink.addEventListener('click', function (e) {         if (dashboardLink) {                  const dashboardLink = document.getElementById('dashboardLink');     document.addEventListener('DOMContentLoaded', function () { <script> ad  �	  =
     $       �  �  q    �  �  9  �  �  T          �  �  �  �  M    �  �  �  ]  Q  -     �
  �
  �
  �
  ^
  P
  E
  >
  =
  <
  ;
  :
  9
  8
  7
  6
  5
  4
  3
  2
  1
  0
  /
  .
  -
  ,
  +
  *
  )
  (
  '
  &
  %
  $
  �	  �	  n	  	  �  �  �  �  |  a  B  �  �  �  P  ;  )      �  �    �  �  �  �  n  /  '  &    �  �  �  �  e  F  '    �  �  �  �  �  �      @php  @endforeach   @endphp       ]);           $selected->profile6           $selected->profile5,           $selected->profile4,           $selected->profile2,           $selected->profile1,           $selected->profile3,       $images = array_merge($images, [       // Collect all profile images into the array   @php @foreach($selecteds as $selected)  @endphp   $images = []; // Initialize an empty array to collect images   $selecteds = App\Models\Selected::inRandomOrder()->take(3)->get();   // Fetch 3 random selected records   @php   <!-- Carousel items -->   </ol>     <li data-target="#carousel" data-slide-to="2"></li>     <li data-target="#carousel" data-slide-to="1"></li>     <li data-target="#carousel" data-slide-to="0" class="active"></li>   <ol class="carousel-indicators">   	<div id="carousel" class="carousel slide carousel-fade" data-ride="carousel">   <div class="banner-container">  <section id="home"> <div id="#top"></div> <!--/.header--> </header>   <!--/.container-->    </div>     <!--/.navbar-->      </nav>       <!--/.navbar-collapse-->        </div>     </ul>     @endif         @endauth         @endif             <li><a href="{{ route('register') }}" class="scroll-link">Register</a></li>         @if (Route::has('regi                                 <a href="{{ route('notifications.markAllRead') }}" id="markAsRead"                                                                                                               {{ $notification->data['action'] }}: {{ $notificatio                                      <a href="{{ $notificat                                               @foreach(auth()->user()->unreadNotificati                          <ul i                          <                      <div id="notificationDropdown" class="notification-dropdown" st                      <!-- Noti                                               <span class="badge" id="notificationCount">{{ auth()->user()->unreadNotificatio                              <i class="fas fa-bell"></i> <!-- Font                           <a href="javascript:void(0)" i                      <div class                      <!--                          @endif     @endif         </li>             <a href="{{ url('/dashboard') }}" class="scroll-link">Dashboard</a>         <li>     @else         </li>             <a href="#" id="dashboardLink" class="scroll-link">Dashboard</a>         <li>     @if ($userStatus === 'pending')     @endphp         $userStatus = auth()->user()->status;     @php @elseif (auth()->user()->user_type === 'rental_owner')     <li><a href="{{ url('/dashboard') }}" class="scroll-link">Dashboard</a></li> @elseif (auth()->user()->user_type === 'tenant')     <li><a href="{{ route('contact.form') }}" class="scroll-link">Dashboard</a></li>        @if (auth()->user()->user_type === 'admin')  	  @auth           @if (Route::has('login'))  		 		@endif 	  <li><a href="#contactUs" class="scroll-link">Contact Us</a></li>          @if (auth()->user()->user_type === 'tenant' || auth()->user()->user_type === 'rental_owner') 	  <li><a href="#team" class="scroll-link">Team</a></li>           <li><a href="#toptenant" class="scroll-link">Top 5</a></li>           <li><a href="#work" class="scroll-link">Highlights Room</a></li>           <li><a href="#aboutUs" class="scroll-link">About Us</a></li>           <li><a href="#location" class="scroll-link">Location</a></li>           <li class="active" id="firstLink"><a href="#home" class="scroll-link">Home</a></li>         <ul class="nav navbar-nav" id="mainNav">       <div id="main-nav" class="collapse navbar-collapse" style>       <!--/.navbar-header--> ad  j   &     h       �  �  �  e  ]  \  �  �  �  7  +  �  �  G  2          �  �  A  :  9    �  u  n  l  a  `  _  Z    �
  �
  �
  �
  V
   
  �	  �	  �	  �	  �	  �	  �	  �	  ~	  k	  N	  5	  	  �  �  �  �  �  a  5    	  �  �  �  �  z  >  �  �  �  �  �  ^  :  '  �  �  z  x  w  N  +    �  �  �  �  �  �  o  .    �  �  k  D    �  �  �  �  a  &  %                                                                                                                            <option value="{{ $hubrental->address }}">             @if($hubrental->status !== 'pending')         @foreach($hubrentals as $hubrental)         </option>             @endif                 List of rental hubs             @elseif (auth()->user()->user_type === 'admin')                 Select your rental hub             @elseif (auth()->user()->user_type === 'rental_owner')                 Select a rental hub             @if (auth()->user()->user_type === 'tenant')         <option selected disabled>     <select id="hubrental-select-dropdown" class="form-control">     <!-- Dropdown for selecting hub rentals --> <div class="dropdown-container">  </style>  }     box-shadow: 0 0 5px rgba(0, 123, 255, 0.5);     outline: none;     border-color: #007bff; #hubrental-select-dropdown:focus { /* Style when the dropdown is focused */  }     overflow: hidden; /* Hide any overflow text */     white-space: nowrap; /* Prevent text from wrapping */     text-overflow: ellipsis; /* Add ellipsis to long options */     padding: 10px; #hubrental-select-dropdown option { /* Style for options in the dropdown */  }     overflow: hidden; /* Hide any overflow text */     white-space: nowrap; /* Prevent the text from wrapping */     text-overflow: ellipsis; /* Add ellipsis when text overflows */     margin-bottom: 20px; /* Add space below the dropdown */     box-shadow: 0 2px 5px rgba(0, 0, 0, 0.1);     color: #333;     background-color: #fff;     border-radius: 4px;     border: 1px solid #ccc;     font-size: 16px;     padding: 6px 12px;     max-width: 420px; /* Set a max-width */     width: 80%; /* Adjust width of the dropdown */ #hubrental-select-dropdown { /* Styling for the dropdown itself */  }     width: 100%; /* Make sure it takes full width for centering */     text-align: center;     align-items: center;     justify-content: center;     display: flex; .dropdown-container { /* Custom style for the dropdown container */ <style>    </div> @endif <h3>Homies Location</h3>   @else   <h3>Add Your Homies Location</h3>    @if (auth()->user()->user_type === 'rental_owner')   <div class="container hero-text2" id="location">  @endphp $tenantprofiles = \App\Models\Tenantprofile::where('user_id', Auth::id())->get(); $hubrentals = \App\Models\Hubrental::all(); $hubrentals = \App\Models\Hubrental::where('user_id', Auth::id())->get(); @php     </div>   	 </div>   <a class="carousel-control right" href="#carousel" data-slide="next">&rsaquo;</a>   <a class="carousel-control left" href="#carousel" data-slide="prev">&lsaquo;</a>   <!-- Carousel controls -->  </div>   <a class="carousel-control right" href="#carousel" data-slide="next">&rsaquo;</a>   <a class="carousel-control left" href="#carousel" data-slide="prev">&lsaquo;</a>   <!-- Carousel controls -->    </div>       @endif           @endforeach               </div>                   <img src="{{ $image }}" alt="banner" style="width: 100%; height: 100%; object-fit: cover;"/>               <div class="item {{ $key === 0 ? 'active' : '' }} fade">           @foreach($images as $key => $image)       @else         <p style="margin: 0; font-size: 30px; color: #333;">No Room Images available.</p> <!-- Message when no images are available -->       @if(empty($images))   <div class="carousel-inner"> <div id="carousel" class="carousel slide" data-ride="carousel"> <!-- Adjust the value as needed -->  @endphp   $images = array_slice($images, 0, 3);   // Limit to a maximum of 3 images   $images = array_filter($images);   // Remove any empty values from the array ad     �     Z       �    l  X  J  C  B  7  6  �  �  B  �  �  l  Q  �  �  �  �  �  �  L  K  0  �  �  r  q  O         �
  �
  �
  �
  n
  
  �	  �	  �	  V	  	  �  �    �  c    �  �  l    �  �  �  �  �  �  W    �  �  �  �  �  �  Q  #  "  �  �  �  �  W  !        �  �  �  z  F      �  �  �  �                                         @if (auth()->user()->user_type === 'rental_owner')              map.setView([userLat, userLng], 13);              var userLng = position.coords.longitude;             var userLat = position.coords.latitude;         navigator.geolocation.getCurrentPosition(function (position) {     if (navigator.geolocation) { function getGeolocation() { // Geolocation function  });     }         selectedHub.marker.openPopup(); // Open popup         map.setView(selectedHub.latlng, 13); // Center the map     if (selectedHub) {      var selectedHub = rentalHubs.find(hub => hub.address === selectedAddress);     // Find the corresponding marker      var selectedAddress = event.target.value; document.getElementById('hubrental-select-dropdown').addEventListener('change', function (event) { // Handle dropdown change event  @endforeach     @endif         });             marker: marker             latlng: [{{ $hubrental->lat }}, {{ $hubrental->lng }}],             address: "{{ $hubrental->address }}",         rentalHubs.push({              `);                 @endauth                     @endif                         @endif                             <a href="/booking-messages/create" class="btn btn-primary">Book Now?</a>                         @else                             <a href="/tenantprofiles" class="btn btn-primary">Book Now?</a>                         @if($tenantprofiles->isEmpty())                     @elseif (auth()->user()->user_type === 'tenant')                         <a href="/selecteds" class="btn btn-primary">View RM</a>                         <a href="/selecteds/create" class="btn btn-primary">Add Room</a>                         <a href="{{route('hubrentals.show',$hubrental->id)}}" class="btn btn-primary">Edit Location</a>                     @if (auth()->user()->user_type === 'rental_owner' && auth()->user()->id === $hubrental->user_id)                 @auth                 Price: P{{ number_format($hubrental->price, 2) }}<br>                 Type: {{ $hubrental->type }}<br>                 {{ $hubrental->address }}<br>                 <b>Owner Name: {{ $hubrental->name }}</b><br>             .bindPopup(`         var marker = L.marker([{{ $hubrental->lat }}, {{ $hubrental->lng }}]).addTo(markersLayer)     @if($hubrental->status !== 'pending') @foreach($hubrentals as $hubrental) // Add markers and populate rental hubs array  var rentalHubs = []; // Array to store rental hubs  var markersLayer = L.featureGroup().addTo(map); // Feature group to store markers  }).addTo(map);     attribution: '&copy; <a href="https://www.openstreetmap.org/copyright">OpenStreetMap</a> contributors' L.tileLayer('https://{s}.tile.openstreetmap.org/{z}/{x}/{y}.png', { // Add OpenStreetMap tiles  var map = L.map('mapid').setView([51.505, -0.09], 13); // Default center // Initialize the map  <script>  <section class="page-section colord" id="mapid" style="height:450px;"> <script src="https://unpkg.com/leaflet-search/dist/leaflet-search.min.js"></script> <!-- Leaflet Search JS --> <link rel="stylesheet" href="https://unpkg.com/leaflet-search/dist/leaflet-search.min.css" /> <!-- Leaflet Search CSS --> <script src="https://unpkg.com/leaflet-control-geocoder/dist/Control.Geocoder.js"></script> <script src="https://unpkg.com/leaflet/dist/leaflet.js"></script> <link rel="stylesheet" href="https://unpkg.com/leaflet-control-geocoder/dist/Control.Geocoder.css" /> <link rel="stylesheet" href="https://unpkg.com/leaflet/dist/leaflet.css" />  </section>  </div>     </select>         @endforeach             @endif                 </option>                     {{ Str::limit($hubrental->name, 40) }} - {{ Str::limit($hubrental->address, 40) }} ad     �     g       �  �  u  =  �  �  ;      �  �  n  >    	  �  �  `  T  G      �  �  �  �  �  �  �  �  �  �  j  .  %    �
  �
  �
  �
  Z
  

  �	  �	  �	  �	  �	  �	  �	  �	  {	  T	  =	  %	    	  �  �  �  �      �  �  �  M  E  D  "    �  �  �  �  d  E  &    �  �  �  �  �  �  �  n  F  >  *    �  �  �  �  ^  )        
  �  �  �        						<div class="col-md-4 col-sm-6">     <div class="row dataTxt">	     </div>  @endif @endforeach     </div>         <img src="{{ $image }}" alt="" width="100%">     <div class="area2 columns feature-media left"> @foreach($images as $image) @else </div>   <p style="color:greenyellow;font-size:20px;">No images room available</p> <div class="col-md-12 text-center"> @if(empty($images)) @endphp   $images = array_slice($images, 0, 1);   // Limit to a maximum of 3 images   $images = array_filter($images);   // Remove any empty values from the array @php  @endforeach   @endphp       ]);           $selected->profile3,           $selected->profile6,           $selected->profile5,           $selected->profile2,           $selected->profile1,           $selected->profile4,       $images = array_merge($images, [       // Collect all profile images into the array   @php @foreach($selecteds as $selected)  @endphp   $images = []; // Initialize an empty array to collect images   $selecteds = App\Models\Selected::inRandomOrder()->take(1)->get();   // Fetch 3 random selected records       @php       </div>         <p>Whether you're looking for comfort or style, our design delivers both, ensuring a space that feels both contemporary and timeless."</p>         <p>"Our spaces are thoughtfully designed with a modern aesthetic and a focus on simplicity and functionality. Each room features clean lines, minimalist decor, and high-quality materials to create a fresh, inviting atmosphere.  </p>         <h3>Clean and Modern Design.</h3>       <div class="area1 columns right">     <div class="row feature design">     </div>       <p>"At Homies, we are dedicated to delivering exceptional experiences. Our journey has been shaped by passion, innovation, and a commitment to excellence. With a focus on quality and customer satisfaction, we continuously strive to meet and exceed expectations."</p>       <h2>About Us</h2>       <!-- Heading -->     <div class="heading text-center">    <div class="container"> <section id="aboutUs">  </script>     });         }             });                 );                     'warning'                     'Your account is still pending. Please wait for approval.',                     'Account Pending',                 Swal.fire(                                  e.preventDefault();             pending.addEventListener('click', function (e) {         if (pending) {                  const pending = document.getElementById('pending');     document.addEventListener('DOMContentLoaded', function () { <script>  </section>  </script>  getGeolocation(); // Center map on user's location  }     }         alert("Geolocation is not supported by your browser.");     } else {         });             alert("Could not get your location. Using default location.");             console.error("Geolocation error:", error.message);         }, function (error) {             @endif                     .openPopup();                     .bindPopup(`You are Here!`)                 L.marker([userLat, userLng]).addTo(map)             @elseif (auth()->user()->user_type === 'tenant')                     .openPopup();                     `)                         @endif                             <a href="{{route('hubrentals.create')}}" class="btn btn-primary" style="height:33px;">Add</a>                         @else                             <a href="#" id="pending" class="btn btn-primary" style="height:33px;">Add</a>                         @if ($userStatus === 'pending')                         Add Your Rental Space<br>                     .bindPopup(`                 L.marker([userLat, userLng]).addTo(map) ad     �     V       �  �  P  D  7  0  
    �  �  Z  4    �  �  �  �  �  �  �  m    �
  �
  �
  �
  o
  0
  �	  �	  �	  |	  Q	  &	  �  �  �  �  �  �  c  6  	  �  �  �  �  q      �  �  �  ]  F  .      
  �  �  �  �  h  �  �  x  Z  =  .  �  �  �  |    �  �  /        �  �  �  �  �  �                             @php   @foreach($selecteds as $selected)      @endphp       $images = []; // Initialize an empty array to collect images       @php       @else           </li>               <p>No Image Room available.</p> <!-- Message when no items are available -->           <li class="item branding" style="width: 100%; text-align: center;background-color:greenyellow;">       @if($selecteds->isEmpty())   <ul class="items list-unstyled clearfix animated fadeInRight showing" data-animation="fadeInRight">   <div class="items-container">       @endphp       $selecteds = App\Models\Selected::inRandomOrder()->take(8)->get();        // Fetch all selected records and randomly select 8           @php         <div id="portfolio">       <div class="col-md-12">     <div class="row">     </div>       <p>"Experience unmatched comfort with a cozy atmosphere and modern decor. This room features a spacious layout, natural lighting, and elegant furnishings, perfect for relaxation and productivity."</p>       <h2>8 Highlights Room Images</h2>     <div class="heading">   <div class="container text-center"> <section id="work" class="page-section page"> </section>    </div> 					</div>         @endif             @endforeach                 </div>                     <img src="{{ $image }}" alt="" width="100%">                 <div class="col-md-4 col-sm-6">             @foreach($images as $image)         @else             </div>                 <p style="color:greenyellow;font-size:20px;">No images room available</p>             <div class="col-md-12 text-center">         @if(empty($images))                   @endphp             $images = array_slice($images, 0, 1);             // Limit to a maximum of 1 image             $images = array_filter($images);             // Remove any empty values from the array             @php                          @endforeach               @endphp                   ]);                       $selected->profile3,                       $selected->profile1,                       $selected->profile4,                       $selected->profile2,                       $selected->profile6,                       $selected->profile5,                   $images = array_merge($images, [                   // Collect all profile images into the array               @php             @foreach($selecteds as $selected)                          @endphp               $images = []; // Initialize an empty array to collect images               $selecteds = App\Models\Selected::inRandomOrder()->take(1)->get();               // Fetch 3 random selected records               @php 							</div> 							<!-- Accordion starts --> 							</ul> 								<li>Our commitment to excellence and attention to detail ensure a seamless experience from start to finish, making us the perfect choice for your living needs."</li> 								<li>we create spaces that truly feel like home.</li> 								<li>and exceptional customer service,</li> 								<li>high-quality amenities,</li> 								<li>With modern designs,</li>                             <ul class="listArrow"> 							<p>"At Homies, we prioritize your comfort, convenience, and satisfaction. </p> 							<h4>Why Choose Us?</h4> 							 						<div class="col-md-4 col-sm-6"> 						 						</div> 							<br>                             <p>Our team works hard to ensure every detail is perfect, delivering exceptional service and a welcoming environment."</p> 							<p>"At Homies, we specialize in creating comfortable, stylish living spaces that cater to your needs. From providing modern, well-designed rooms to offering a seamless rental experience, we are dedicated to making your stay feel like home.  </p> 							<h4>What We Do?</h4> ad  =        m       �  �  {  X  5    �  �  �  �  �  �  �  i  B    �  �  �  �  S    �  �  p  (    �  �  �  �  �  �  �  �  �  �  �  u  G  -    �
  �
  y
  =
  2
  
  �	  �	  �	  �	  :	  	  �  �  �  �  d  ?  >    �  �  u  D  
  �  �  �  �  �  �  Q  C  8  7  6    �  �  �  +  �  �  �  �  �  �  �  �  �  L  1      �  �  �  �  �  e    �  �  �  \  4                                                                                       {{ $index + 1 }}.                  <li class="plan-price">             @foreach ($bookingmessages as $index => $bookingmessage)         @else             <li class="plan-price">No Booking yet.</li>         @if ($bookingmessages->isEmpty())         <!-- Show booking list for all user types (tenant, rental_owner, admin) -->         <li class="plan-name">Top Book List</li>     <ul class="plan plan2 featured"> <div class="col-lg-3 col-md-3 col-sm-6 col-xs-12">  @endphp     ->get();     ->take(5)     ->orderBy('count', 'desc')     ->groupBy('sender_id') $bookingmessages = \App\Models\BookingMessage::selectRaw('sender_id, COUNT(*) as count') @php   </div>       </ul>         </li>         @endif             @endforeach                 {{-- ({{ $tenant->login_count }}) --}}                 <li class="plan-price">{{ $index + 1 }}. <strong>{{ $tenant->name }}</strong></li>             @foreach ($tenants as $index => $tenant)         @else             <li class="plan-price">No tenants registered yet.</li>         @if ($tenants->isEmpty())       @endif     @endguest         <li class="plan-name">Top Name List</li>     @guest @else     @endif         <li class="plan-name">Top Name List</li>     @else         <li class="plan-name">Top Name List</li>     @elseif(auth()->user()->user_type === 'rental_owner')         <li class="plan-name">Top Name List</li>     @if (auth()->user()->user_type === 'tenant') @elseif (auth()->check())     <li class="plan-name"><a href="{{ route('register') }}">Register?</a></li> @if (!auth()->check() && $registeredCount < 5)      <ul class="plan plan2 featured"> <div class="col-lg-3 col-md-3 col-sm-6 col-xs-12"> 		 @endphp 	$registeredCount = \App\Models\User::count(); // Count all registered users 	->get(); // Get top 5 tenants         ->take(5) // Limit to top 5 tenants         ->orderBy('login_count', 'desc') // Sort by login_count in descending order     $tenants = App\Models\User::where('user_type', 'tenant')  @php       </div>       <div class="col-lg-3 col-md-3 col-sm-6 col-xs-12">     <div class="row flat">     </div>       <p>Book now and get access to our top 5 bookings.</p>       <p>Register now  and get access to our top 5 visitors.</p>       <h2>The Top 5 Tenant Visitors And Booking</h2>       <!-- Heading -->     <div class="heading text-center">    <div class="container"> <section id="toptenant" class="page-section"> </section>   </div>     </div>       </div>         </div>        </div>      </ul>      @endif        @endforeach           </li>           </figure>               </figcaption>                   <a href="{{ $image }}" class="fancybox">View more</a>                   <h2>Trends</h2>               <figcaption>               <img src="{{ $image }}" alt="Image" style="width: 100%; height: 200px; object-fit: cover;"/>           <figure class="effect-bubba" style="margin: 0;">       <li class="item branding" style="display: inline-block; width: 25%; box-sizing: border-box; padding: 0;">   @foreach($images as $image)      @endphp       $images = array_slice($images, 0, 8);       // Limit to a maximum of 8 images       $images = array_filter($images);       // Remove any empty values from the array   @php      @endforeach       @endphp           ]);               $selected->profile6               $selected->profile5,               $selected->profile4,               $selected->profile3,               $selected->profile2,               $selected->profile1,           $images = array_merge($images, [           // Collect all profile images into the array ad  4   �     X       �  y  a  R  H  A  @    �  �  �  �  �  �  l  R  +       �  �  ^  ?  '  �  �  �  �  ]  >  �  �  �  h  F    �
  
  
  �	  �	  �	  |	  U	  /	  	  �  �  b  @    w  f  W  $    �  �  �  n    �  �  �  Y  �  �  �  s  T  )    �  �  U  1    �  �      �  �  �  �  �  �  �  �                                                       </section>   <!--/.container-->    </div>     </div>       </div>         </div>           </div>             <div class="team-socials"> <a href="https://www.facebook.com/hartjadefranz.gallego" target="_blank"><i class="fa fa-facebook"></i></a></div>             <span class="pos">The Documentator</span>             <!-- Designation -->              <h4>Hartjade Franz Gallego </h4>             <!-- Member Details -->               <img class="img-responsive" src="10.jpg" alt=""  style="height:150px;width:200px"> </div>               <!-- Image  -->              <div class="member-img">              <!-- Image Hover Block -->           <div class="team-member pDark">            <!-- Team Member -->         <div class="col-md-3 col-sm-6 col-xs-12">          </div>           </div>             <div class="team-socials"> <a href="https://www.facebook.com/princejoao.caya" target="_blank"><i class="fa fa-facebook"></i></a></div>             <span class="pos">The System Analys</span>             <!-- Designation -->              <h4>Esteve Mark Salamanca Caya</h4>             <!-- Member Details -->               <img class="img-responsive" src="11.jpg" alt=""  style="height:150px;width:200px"> </div>               <!-- Image  -->              <div class="member-img">              <!-- Image Hover Block -->           <div class="team-member pDark">            <!-- Team Member -->         <div class="col-md-3 col-sm-6 col-xs-12">          </div>           </div>             <div class="team-socials"> <a href="https://github.com/germanybasillo" target="_blank"><i class="fa fa-github"></i></a></div>             <span class="pos">The Programmer / Designer</span>             <!-- Designation -->              <h4>Germany Lungay</h4>             <!-- Member Details -->               <img class="img-responsive" src="9.jpg" alt="" style="height:150px;width:200px"> </div>               <!-- Image  -->              <div class="member-img">              <!-- Image Hover Block -->           <div class="team-member pDark">            <!-- Team Member -->         <div class="col-md-3 col-sm-6 col-xs-12">          </div>           </div>             <div class="team-socials"> <a href="https://www.facebook.com/Miharbe.diangca" target="_blank"><i class="fa fa-facebook"></i><a href="https://github.com/ediangca" target="_blank"><i class="fa fa-github"></i></a> </div> 			    </div>             <span class="pos">Our Teacher Adviser</span>             <!-- Designation -->  		      	<h4>Mr. Ebrahim Diangca</h4>             <div class="team-title">             <!-- Member Details -->               <img class="img-responsive" src="8.jpg" alt=""  style="height:150px;width:200px"> </div>               <!-- Image  -->              <div class="member-img">              <!-- Image Hover Block -->           <div class="team-member pDark">            <!-- Team Member -->         <div class="col-md-3 col-sm-6 col-xs-12">        <div class="row">     <div class="team-content">     <!-- Team Member's Details -->     </div>       <p>Driven by passion and dedication, our team is here to make a difference in every project we undertake.</p>       <h2>Team</h2>       <!-- Heading -->     <div class="heading text-center">    <div class="container"> <section id="team" class="page-section"> </section>   </div>     </div>       </div>       <div class="col-lg-3 col-md-3 col-sm-6 col-xs-12">       </div>       <div class="col-lg-3 col-md-3 col-sm-6 col-xs-12">  </div>     </ul>         @endif             @endforeach                 </li>                     <strong>{{ $bookingmessage->sender->name }}</strong> ({{ $bookingmessage->count }} bookings) ad     }     Q       �  �  r  V  :  "  �  �  �  �  �  �  �  �  �  G  7    �  �  �  �  w  D  N
  9
  
  �	  �  �  w  I  8  *  )  (    �  �  �  E  �  �  �  �  �  v  ^  ?    �  �  �  �  �  �  2  �  �  �  g  	  �  �  �  c  ;  +  �  �  �  �  �  �  \  +    �  �  �  }  |                                       .then(data => {         .then(response => response.json()) // Assuming your controller returns JSON         })             body: formData             method: "POST",         fetch("{{ route('contact.submit') }}", {         // Use AJAX to submit the form          var formData = new FormData(this);         // Create a FormData object to handle the form data          }             return; // Stop the form from submitting             });                 confirmButtonText: 'OK'                 text: 'You can only submit the form once every 24 hours.',                 title: 'Oops...',                 icon: 'warning',             Swal.fire({         if (lastSubmissionTime && (currentTime - lastSubmissionTime < 24 * 60 * 60 * 1000)) {         // If the last submission was within the last 24 hours          const currentTime = new Date().getTime();         const lastSubmissionTime = localStorage.getItem('lastSubmissionTime_' + userId);         // Check the last submission time for the specific user in localStorage          }             return;             });                 confirmButtonText: 'OK'                 text: 'You need to be logged in to submit the form.',                 title: 'Error',                 icon: 'error',             Swal.fire({         if (!userId) {         // Check if the user is logged in          const userId = {{ Auth::check() ? Auth::id() : 'null' }};           e.preventDefault(); // Prevent the form from submitting normally     document.getElementById('contactfrm').addEventListener('submit', function(e) {     // Listen for the form submission <script> <script src="https://cdn.jsdelivr.net/npm/sweetalert2@11"></script> <!-- Include SweetAlert2 -->         </form>           </div>               <div class="result mt-3"></div>               <button name="submit" type="submit" class="btn btn-lg btn-primary">Submit</button>               </div>                   <textarea name="comment" class="form-control" id="comments" cols="3" rows="5" placeholder="Enter your message…" required minlength="10" title="Please enter your message (at least 10 characters)" required></textarea>                   <label for="comments">Comments</label>               <div class="form-group">               </div>                   <input type="email" class="form-control" name="email" id="email" value="{{ Auth::user()->email ?? null }}"   {{ Auth::check() ? 'readonly' : '' }}  required  placeholder="Enter Email" title="Please enter a valid email address">                   <label for="email">Email</label>               <div class="form-group">               </div>                   <input type="text" class="form-control" name="name" id="name" value="{{ Auth::user()->name ?? null }}"   {{ Auth::check() ? 'readonly' : '' }}  required minlength="2" placeholder="Enter name" title="Please enter your name (at least 2 characters)">                   <label for="name">Name</label>               <div class="form-group">           <div class="col-sm-12">           @csrf         <form method="post" action="{{ route('contact.submit') }}" id="contactfrm" role="form" novalidate>         <div class="row mrgn30">       </div>         </div>           <p>"We’re here to help! Reach out to us with any questions, and our team will be happy to assist you. Whether you need more information or have specific requests, feel free to get in touch."</p>           <h2>Contact Us</h2>           <!-- Heading -->         <div class="heading text-center">        <div class="row">     <div class="container">   <div class="parlex-back"> <section id="contactUs" class="contact-parlex">  @if (auth()->user()->user_type === 'tenant' || auth()->user()->user_type === 'rental_owner') ad      �     f       �  �  �  p  G  �  �  }    �  �  A  -    �  �  �  {  &  �  �  �  �  �  �  o  P  .  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  }
  r
  Z
  Q
  F
  ?
  )
  
  �	  �	  �	  �	  L	  	  �  �  �  x  c  Z  O      �  T    �  \  �  �  u  @  �  �  o  f  (    �  �  �  x  j  D  .    �  �  �  �  �  �  �  �  T  -    �  �                showNoInternetMessage();           // If no internet connection, show a message       if (!navigator.onLine) {   function checkInternetConnection() {   // Function to check if the browser is offline <script>    </script>   });       @endif           });               text: '{{ session('swal:login') }}',               title: 'Success',               icon: 'success',           Swal.fire({       @elseif (session('swal:login'))           });               text: '{{ session('swal:register') }}',               title: 'Success',               icon: 'success',           Swal.fire({       @if (session('swal:register'))   document.addEventListener('DOMContentLoaded', function () { <script> <script src="https://cdn.jsdelivr.net/npm/sweetalert2@11"></script> <script src="landingpage/js/owl-carousel/owl.carousel.js"></script> <script src="landingpage/js/custom.js" type="text/javascript"></script>  <script src="landingpage/js/waypoints.js"></script>  <script src="landingpage/js/jquery.fittext.js"></script>  <script src="landingpage/js/jquery.nav.js" type="text/javascript"></script>  <script src="landingpage/js/fancybox/jquery.fancybox.pack.js" type="text/javascript"></script>  <script src="landingpage/js/jquery.isotope.min.js" type="text/javascript"></script>  <script src="landingpage/js/bootstrap.min.js" type="text/javascript"></script>  <script src="landingpage/js/jquery-1.8.2.min.js" type="text/javascript"></script>  <script src="landingpage/js/modernizr-latest.js"></script>  <!--[if lte IE 8]><script src="//ajax.googleapis.com/ajax/libs/jquery/1.11.0/jquery.min.js"></script><![endif]-->   <a href="#top" class="topHome"><i class="fa fa-chevron-up fa-2x"></i></a>  </section>   </div>     <!-- / .row -->      </div>       </script>         });           document.getElementById('copyright').innerHTML = `Copyright ${year} | All Rights Reserved -- Homies - Capstone2`;           const year = new Date().getFullYear();         document.addEventListener("DOMContentLoaded", function() {       <script>       <div class="col-sm-12 text-center" id="copyright"></div>     <div class="row">   <div class="container"> <section class="copyright"> <!--/.page-section--> @endif </section>   </div>     <!--/.container-->      </div>     </div>          </script>     });         });             });                 confirmButtonText: 'OK'                 text: 'An error occurred while sending your message.',                 title: 'Oops...',                 icon: 'error',             Swal.fire({             console.error('Error:', error);         .catch(error => {         })             }                 });                     confirmButtonText: 'OK'                     text: data.message || 'Something went wrong, please try again.',                     title: 'Oops...',                     icon: 'error',                 Swal.fire({                 // Show error message if not successful             } else {                 });                     document.getElementById('contactfrm').reset();                     // Optionally, reset the form                     localStorage.setItem('lastSubmissionTime_' + userId, currentTime);                     // Save the current time in localStorage to prevent another submission in the next 24 hours                 }).then(() => {                     confirmButtonText: 'OK'                     text: data.message || 'Your message has been successfully submitted. Wait for the admin to contact you!',                     title: 'Thank you!',                     icon: 'success',                 Swal.fire({                 // Show SweetAlert2 on success             if (data.success) { 